// cpu.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module cpu (
		output wire [15:0] apple_o_export,      //      apple_o.export
		input  wire        clk_clk,             //          clk.clk
		output wire [15:0] erace_o_export,      //      erace_o.export
		input  wire [1:0]  movement_i_export,   //   movement_i.export
		input  wire        rst_n_i_export,      //      rst_n_i.export
		output wire [7:0]  score_o_export,      //      score_o.export
		output wire [15:0] snake_head_o_export  // snake_head_o.export
	);

	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [15:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [15:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;           // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;             // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;              // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;           // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;            // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_rst_n_i_s1_readdata;                      // rst_n_i:readdata -> mm_interconnect_0:rst_n_i_s1_readdata
	wire   [1:0] mm_interconnect_0_rst_n_i_s1_address;                       // mm_interconnect_0:rst_n_i_s1_address -> rst_n_i:address
	wire  [31:0] mm_interconnect_0_movement_i_s1_readdata;                   // movement_i:readdata -> mm_interconnect_0:movement_i_s1_readdata
	wire   [1:0] mm_interconnect_0_movement_i_s1_address;                    // mm_interconnect_0:movement_i_s1_address -> movement_i:address
	wire         mm_interconnect_0_apple_o_s1_chipselect;                    // mm_interconnect_0:apple_o_s1_chipselect -> apple_o:chipselect
	wire  [31:0] mm_interconnect_0_apple_o_s1_readdata;                      // apple_o:readdata -> mm_interconnect_0:apple_o_s1_readdata
	wire   [1:0] mm_interconnect_0_apple_o_s1_address;                       // mm_interconnect_0:apple_o_s1_address -> apple_o:address
	wire         mm_interconnect_0_apple_o_s1_write;                         // mm_interconnect_0:apple_o_s1_write -> apple_o:write_n
	wire  [31:0] mm_interconnect_0_apple_o_s1_writedata;                     // mm_interconnect_0:apple_o_s1_writedata -> apple_o:writedata
	wire         mm_interconnect_0_snake_head_o_s1_chipselect;               // mm_interconnect_0:snake_head_o_s1_chipselect -> snake_head_o:chipselect
	wire  [31:0] mm_interconnect_0_snake_head_o_s1_readdata;                 // snake_head_o:readdata -> mm_interconnect_0:snake_head_o_s1_readdata
	wire   [1:0] mm_interconnect_0_snake_head_o_s1_address;                  // mm_interconnect_0:snake_head_o_s1_address -> snake_head_o:address
	wire         mm_interconnect_0_snake_head_o_s1_write;                    // mm_interconnect_0:snake_head_o_s1_write -> snake_head_o:write_n
	wire  [31:0] mm_interconnect_0_snake_head_o_s1_writedata;                // mm_interconnect_0:snake_head_o_s1_writedata -> snake_head_o:writedata
	wire         mm_interconnect_0_erace_o_s1_chipselect;                    // mm_interconnect_0:erace_o_s1_chipselect -> erace_o:chipselect
	wire  [31:0] mm_interconnect_0_erace_o_s1_readdata;                      // erace_o:readdata -> mm_interconnect_0:erace_o_s1_readdata
	wire   [1:0] mm_interconnect_0_erace_o_s1_address;                       // mm_interconnect_0:erace_o_s1_address -> erace_o:address
	wire         mm_interconnect_0_erace_o_s1_write;                         // mm_interconnect_0:erace_o_s1_write -> erace_o:write_n
	wire  [31:0] mm_interconnect_0_erace_o_s1_writedata;                     // mm_interconnect_0:erace_o_s1_writedata -> erace_o:writedata
	wire         mm_interconnect_0_score_o_s1_chipselect;                    // mm_interconnect_0:score_o_s1_chipselect -> score_o:chipselect
	wire  [31:0] mm_interconnect_0_score_o_s1_readdata;                      // score_o:readdata -> mm_interconnect_0:score_o_s1_readdata
	wire   [1:0] mm_interconnect_0_score_o_s1_address;                       // mm_interconnect_0:score_o_s1_address -> score_o:address
	wire         mm_interconnect_0_score_o_s1_write;                         // mm_interconnect_0:score_o_s1_write -> score_o:write_n
	wire  [31:0] mm_interconnect_0_score_o_s1_writedata;                     // mm_interconnect_0:score_o_s1_writedata -> score_o:writedata
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [apple_o:reset_n, erace_o:reset_n, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, movement_i:reset_n, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_n_i:reset_n, rst_translator:in_reset, score_o:reset_n, snake_head_o:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	cpu_apple_o apple_o (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_apple_o_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_apple_o_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_apple_o_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_apple_o_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_apple_o_s1_readdata),   //                    .readdata
		.out_port   (apple_o_export)                           // external_connection.export
	);

	cpu_apple_o erace_o (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_erace_o_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_erace_o_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_erace_o_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_erace_o_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_erace_o_s1_readdata),   //                    .readdata
		.out_port   (erace_o_export)                           // external_connection.export
	);

	cpu_movement_i movement_i (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_movement_i_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_movement_i_s1_readdata), //                    .readdata
		.in_port  (movement_i_export)                         // external_connection.export
	);

	cpu_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	cpu_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	cpu_rst_n_i rst_n_i (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_rst_n_i_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_rst_n_i_s1_readdata), //                    .readdata
		.in_port  (rst_n_i_export)                         // external_connection.export
	);

	cpu_score_o score_o (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_score_o_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_score_o_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_score_o_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_score_o_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_score_o_s1_readdata),   //                    .readdata
		.out_port   (score_o_export)                           // external_connection.export
	);

	cpu_apple_o snake_head_o (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_snake_head_o_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_snake_head_o_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_snake_head_o_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_snake_head_o_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_snake_head_o_s1_readdata),   //                    .readdata
		.out_port   (snake_head_o_export)                           // external_connection.export
	);

	cpu_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                    //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.apple_o_s1_address                             (mm_interconnect_0_apple_o_s1_address),                       //                               apple_o_s1.address
		.apple_o_s1_write                               (mm_interconnect_0_apple_o_s1_write),                         //                                         .write
		.apple_o_s1_readdata                            (mm_interconnect_0_apple_o_s1_readdata),                      //                                         .readdata
		.apple_o_s1_writedata                           (mm_interconnect_0_apple_o_s1_writedata),                     //                                         .writedata
		.apple_o_s1_chipselect                          (mm_interconnect_0_apple_o_s1_chipselect),                    //                                         .chipselect
		.erace_o_s1_address                             (mm_interconnect_0_erace_o_s1_address),                       //                               erace_o_s1.address
		.erace_o_s1_write                               (mm_interconnect_0_erace_o_s1_write),                         //                                         .write
		.erace_o_s1_readdata                            (mm_interconnect_0_erace_o_s1_readdata),                      //                                         .readdata
		.erace_o_s1_writedata                           (mm_interconnect_0_erace_o_s1_writedata),                     //                                         .writedata
		.erace_o_s1_chipselect                          (mm_interconnect_0_erace_o_s1_chipselect),                    //                                         .chipselect
		.movement_i_s1_address                          (mm_interconnect_0_movement_i_s1_address),                    //                            movement_i_s1.address
		.movement_i_s1_readdata                         (mm_interconnect_0_movement_i_s1_readdata),                   //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),              //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                         .clken
		.rst_n_i_s1_address                             (mm_interconnect_0_rst_n_i_s1_address),                       //                               rst_n_i_s1.address
		.rst_n_i_s1_readdata                            (mm_interconnect_0_rst_n_i_s1_readdata),                      //                                         .readdata
		.score_o_s1_address                             (mm_interconnect_0_score_o_s1_address),                       //                               score_o_s1.address
		.score_o_s1_write                               (mm_interconnect_0_score_o_s1_write),                         //                                         .write
		.score_o_s1_readdata                            (mm_interconnect_0_score_o_s1_readdata),                      //                                         .readdata
		.score_o_s1_writedata                           (mm_interconnect_0_score_o_s1_writedata),                     //                                         .writedata
		.score_o_s1_chipselect                          (mm_interconnect_0_score_o_s1_chipselect),                    //                                         .chipselect
		.snake_head_o_s1_address                        (mm_interconnect_0_snake_head_o_s1_address),                  //                          snake_head_o_s1.address
		.snake_head_o_s1_write                          (mm_interconnect_0_snake_head_o_s1_write),                    //                                         .write
		.snake_head_o_s1_readdata                       (mm_interconnect_0_snake_head_o_s1_readdata),                 //                                         .readdata
		.snake_head_o_s1_writedata                      (mm_interconnect_0_snake_head_o_s1_writedata),                //                                         .writedata
		.snake_head_o_s1_chipselect                     (mm_interconnect_0_snake_head_o_s1_chipselect)                //                                         .chipselect
	);

	cpu_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
